
class clk_rst_uvc extends uvm_env;
	

	
	`uvm_component_utils(clk_rst_uvc);

	function new(string name = "clk_rst_uvc", uvm_component parent);
		super.new(name, parent);
	endfunction

	
endclass
