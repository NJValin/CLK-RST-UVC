`default_nettype none

interface clk_rst_if (
		input logic clk,
		input logic clkb
	);

	clk_rst_cfg cfg;
	
endinterface
